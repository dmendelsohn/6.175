// The contents of this file has been moved to ProcTypes.bsv (I think...)
